module ex7_top(
KEY,
HEX0,
HEX1
);

	input [3:0] KEY;
	output [6:0] HEX0, HEX1;
	
	wire [6:0] data_out;
	
	LFSR_7 LFSR(data_out, ~KEY[3]);
	
	hex_to_7seg SEG0(HEX0, data_out[3:0]);
	hex_to_7seg SEG1(HEX1, {1'b0, data_out[6:4]});
	
endmodule
